module Gates(
    input in1,in2;
    output out
);
    //assign out=in1;-------->a wire
    //assign out=1'b0;------>VSS(电源负极)GND(接地)
    //assign out=in1&in2---->AND(与门)
endmodule