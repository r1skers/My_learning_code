module Gates(
    input in1,in2;
    output out
);
    //assign out=in1;-------->a wire
    //assign out=1'b0;------>VSS(电源负极)GND(接地)
    //assign out=in1&in2;---->AND(与门)
    //assign out=in1|in2;---->OR(或门)
    //assign out=~in1;------->INVERTER(非门)
    //assign out=~(in1|in2);->NOR(或非门)
    //assign out=in1^in2;---->XOR(异或门)
    //assign out=~(in1&in2);->NAND(与非门)
    //assign out=~(in1^in2);->XNOR(同或门)
endmodule
