module Gates();